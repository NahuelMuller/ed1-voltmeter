-------------------------------------------------
-- Memoria	(rom_char)
--
-- Descripcion: Memoria de caracteres
-- Entradas:	Selectores fila y columna
-- Salidas:		Bit pixel
--
-- Autor:		Nahuel Müller
-------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity rom_char is
	port(
		fila: in integer range 0 to 103; 
		columna: in integer range 0 to 7;
		mem_out: out std_logic
	);
end entity;

architecture rom_char_arq of rom_char is

	type mem_104x8 is array (0 to 103, 0 to 7) of std_logic;

	constant char_mem: mem_104x8:= (
								('0','1','1','1','1','1','1','0'),	-- Caracter 0
								('0','1','0','0','0','1','1','0'),
								('0','1','0','0','1','0','1','0'),
								('0','1','0','0','0','0','1','0'),
								('0','1','0','1','0','0','1','0'),
								('0','1','1','0','0','0','1','0'),
								('0','1','1','1','1','1','1','0'),
								('0','0','0','0','0','0','0','0'),
								
								('0','0','0','0','1','0','0','0'),	-- Caracter 1
								('0','0','0','1','1','0','0','0'),
								('0','0','1','0','1','0','0','0'),
								('0','0','0','0','1','0','0','0'),
								('0','0','0','0','1','0','0','0'),
								('0','0','0','0','1','0','0','0'),
								('0','0','1','1','1','1','0','0'),
								('0','0','0','0','0','0','0','0'),
								
								('0','0','1','1','1','1','0','0'),	-- Caracter 2
								('0','1','0','0','0','0','1','0'),
								('0','0','0','0','0','1','0','0'),
								('0','0','0','0','1','0','0','0'),
								('0','0','0','1','0','0','0','0'),
								('0','0','1','0','0','0','0','0'),
								('0','1','1','1','1','1','1','0'),
								('0','0','0','0','0','0','0','0'),
								
								('0','0','1','1','1','1','0','0'),	-- Caracter 3
								('0','1','0','0','0','0','1','0'),
								('0','0','0','0','0','0','1','0'),
								('0','0','0','1','1','1','0','0'),
								('0','0','0','0','0','0','1','0'),
								('0','1','0','0','0','0','1','0'),
								('0','0','1','1','1','1','0','0'),
								('0','0','0','0','0','0','0','0'),
								
								('0','0','0','0','1','1','0','0'),	-- Caracter 4
								('0','0','0','1','0','1','0','0'),
								('0','0','1','0','0','1','0','0'),
								('0','1','0','0','0','1','0','0'),
								('0','1','1','1','1','1','1','0'),
								('0','0','0','0','0','1','0','0'),
								('0','0','0','0','0','1','0','0'),
								('0','0','0','0','0','0','0','0'),
								
								('0','1','1','1','1','1','1','0'),	-- Caracter 5
								('0','1','0','0','0','0','0','0'),
								('0','1','0','0','0','0','0','0'),
								('0','0','1','1','1','1','0','0'),
								('0','0','0','0','0','0','1','0'),
								('0','1','0','0','0','0','1','0'),
								('0','0','1','1','1','1','0','0'),
								('0','0','0','0','0','0','0','0'),
								
								('0','0','1','1','1','1','0','0'),	-- Caracter 6
								('0','1','0','0','0','0','1','0'),
								('0','1','0','0','0','0','0','0'),
								('0','1','1','1','1','1','0','0'),
								('0','1','0','0','0','0','1','0'),
								('0','1','0','0','0','0','1','0'),
								('0','0','1','1','1','1','0','0'),
								('0','0','0','0','0','0','0','0'),
								
								('0','1','1','1','1','1','1','0'),	-- Caracter 7
								('0','1','0','0','0','0','1','0'),
								('0','0','0','0','0','1','1','0'),
								('0','0','0','0','1','1','0','0'),
								('0','0','0','0','1','0','0','0'),
								('0','0','0','1','0','0','0','0'),
								('0','0','0','1','0','0','0','0'),
								('0','0','0','0','0','0','0','0'),
								
								('0','0','1','1','1','1','0','0'),	-- Caracter 8
								('0','1','0','0','0','0','1','0'),
								('0','1','0','0','0','0','1','0'),
								('0','0','1','1','1','1','0','0'),
								('0','1','0','0','0','0','1','0'),
								('0','1','0','0','0','0','1','0'),
								('0','0','1','1','1','1','0','0'),
								('0','0','0','0','0','0','0','0'),
								
								('0','0','1','1','1','1','0','0'),	-- Caracter 9
								('0','1','0','0','0','0','1','0'),
								('0','1','0','0','0','0','1','0'),
								('0','0','1','1','1','1','1','0'),
								('0','0','0','0','0','0','1','0'),
								('0','1','0','0','0','0','1','0'),
								('0','0','1','1','1','1','0','0'),
								('0','0','0','0','0','0','0','0'),
								
								('0','0','0','0','0','0','0','0'),	-- Caracter punto decimal
								('0','0','0','0','0','0','0','0'),
								('0','0','0','0','0','0','0','0'),
								('0','0','0','0','0','0','0','0'),
								('0','0','0','0','0','0','0','0'),
								('0','0','0','1','1','0','0','0'),
								('0','0','0','1','1','0','0','0'),
								('0','0','0','0','0','0','0','0'),
								
								('0','1','0','0','0','0','1','0'),	-- Caracter V
								('0','1','0','0','0','0','1','0'),
								('0','1','0','0','0','0','1','0'),
								('0','1','0','0','0','0','1','0'),
								('0','0','1','0','0','1','0','0'),
								('0','0','0','1','1','0','0','0'),
								('0','0','0','1','1','0','0','0'),
								('0','0','0','0','0','0','0','0'),
								
								('0','0','0','0','0','0','0','0'),	-- Caracter vacio
								('0','0','0','0','0','0','0','0'),
								('0','0','0','0','0','0','0','0'),
								('0','0','0','0','0','0','0','0'),
								('0','0','0','0','0','0','0','0'),
								('0','0','0','0','0','0','0','0'),
								('0','0','0','0','0','0','0','0'),
								('0','0','0','0','0','0','0','0')
								);
begin

	mem_out <= char_mem(fila, columna);

end architecture;